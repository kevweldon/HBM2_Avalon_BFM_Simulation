// ed_sim.v

// Generated using ACDS version 22.4 94

`timescale 1 ps / 1 ps
module ed_sim (
		output wire  sim_checker_traffic_gen_pass,         //        sim_checker.traffic_gen_pass
		output wire  sim_checker_traffic_gen_fail,         //                   .traffic_gen_fail
		output wire  sim_checker_traffic_gen_timeout,      //                   .traffic_gen_timeout
		output wire  cal_status_checker_local_cal_success, // cal_status_checker.local_cal_success
		output wire  cal_status_checker_local_cal_fail     //                   .local_cal_fail
	);

	wire          tg0_0_ctrl_amm_waitrequest;                                             // hbm_0_example_design:ctrl_amm_0_0_waitrequest_n -> tg0_0:amm_ready
	wire  [255:0] tg0_0_ctrl_amm_readdata;                                                // hbm_0_example_design:ctrl_amm_0_0_readdata -> tg0_0:amm_readdata
	wire          tg0_0_ctrl_amm_read;                                                    // tg0_0:amm_read -> hbm_0_example_design:ctrl_amm_0_0_read
	wire   [28:0] tg0_0_ctrl_amm_address;                                                 // tg0_0:amm_address -> hbm_0_example_design:ctrl_amm_0_0_address
	wire   [31:0] tg0_0_ctrl_amm_byteenable;                                              // tg0_0:amm_byteenable -> hbm_0_example_design:ctrl_amm_0_0_byteenable
	wire          tg0_0_ctrl_amm_readdatavalid;                                           // hbm_0_example_design:ctrl_amm_0_0_readdatavalid -> tg0_0:amm_readdatavalid
	wire          tg0_0_ctrl_amm_write;                                                   // tg0_0:amm_write -> hbm_0_example_design:ctrl_amm_0_0_write
	wire  [255:0] tg0_0_ctrl_amm_writedata;                                               // tg0_0:amm_writedata -> hbm_0_example_design:ctrl_amm_0_0_writedata
	wire    [6:0] tg0_0_ctrl_amm_burstcount;                                              // tg0_0:amm_burstcount -> hbm_0_example_design:ctrl_amm_0_0_burstcount
	wire          tg0_1_ctrl_amm_waitrequest;                                             // hbm_0_example_design:ctrl_amm_0_1_waitrequest_n -> tg0_1:amm_ready
	wire  [255:0] tg0_1_ctrl_amm_readdata;                                                // hbm_0_example_design:ctrl_amm_0_1_readdata -> tg0_1:amm_readdata
	wire          tg0_1_ctrl_amm_read;                                                    // tg0_1:amm_read -> hbm_0_example_design:ctrl_amm_0_1_read
	wire   [28:0] tg0_1_ctrl_amm_address;                                                 // tg0_1:amm_address -> hbm_0_example_design:ctrl_amm_0_1_address
	wire   [31:0] tg0_1_ctrl_amm_byteenable;                                              // tg0_1:amm_byteenable -> hbm_0_example_design:ctrl_amm_0_1_byteenable
	wire          tg0_1_ctrl_amm_readdatavalid;                                           // hbm_0_example_design:ctrl_amm_0_1_readdatavalid -> tg0_1:amm_readdatavalid
	wire          tg0_1_ctrl_amm_write;                                                   // tg0_1:amm_write -> hbm_0_example_design:ctrl_amm_0_1_write
	wire  [255:0] tg0_1_ctrl_amm_writedata;                                               // tg0_1:amm_writedata -> hbm_0_example_design:ctrl_amm_0_1_writedata
	wire    [6:0] tg0_1_ctrl_amm_burstcount;                                              // tg0_1:amm_burstcount -> hbm_0_example_design:ctrl_amm_0_1_burstcount
	wire          ref_clk_source_clk_clk;                                                 // ref_clk_source:clk -> [global_reset_n_source:clk, hbm_0_example_design:pll_ref_clk, hbm_only_reset_source:clk]
	wire          core_clk_source_clk_clk;                                                // core_clk_source:clk -> core_clk_iopll:refclk
	wire          core_clk_iopll_outclk0_clk;                                             // core_clk_iopll:outclk_0 -> hbm_0_example_design:ext_core_clk
	wire          hbm_0_example_design_wmc_clk_0_clk;                                     // hbm_0_example_design:wmc_clk_0_clk -> [tg0_0:wmc_clk_in, tg0_1:wmc_clk_in]
	wire    [1:0] tg0_0_apb_ur_pstrb;                                                     // tg0_0:ur_pstrb -> hbm_0_example_design:apb_0_ur_pstrb
	wire   [15:0] tg0_0_apb_ur_pwdata;                                                    // tg0_0:ur_pwdata -> hbm_0_example_design:apb_0_ur_pwdata
	wire          tg0_0_apb_ur_penable;                                                   // tg0_0:ur_penable -> hbm_0_example_design:apb_0_ur_penable
	wire   [15:0] tg0_0_apb_ur_paddr;                                                     // tg0_0:ur_paddr -> hbm_0_example_design:apb_0_ur_paddr
	wire          tg0_0_apb_ur_psel;                                                      // tg0_0:ur_psel -> hbm_0_example_design:apb_0_ur_psel
	wire          tg0_0_apb_ur_pwrite;                                                    // tg0_0:ur_pwrite -> hbm_0_example_design:apb_0_ur_pwrite
	wire          hbm_0_example_design_apb_0_ur_prready;                                  // hbm_0_example_design:apb_0_ur_prready -> tg0_0:ur_prready
	wire   [15:0] hbm_0_example_design_apb_0_ur_prdata;                                   // hbm_0_example_design:apb_0_ur_prdata -> tg0_0:ur_prdata
	wire          hbm_0_example_design_ctrl_ecc_readdataerror_0_0_ctrl_ecc_readdataerror; // hbm_0_example_design:ctrl_ecc_readdataerror_0_0_ctrl_ecc_readdataerror -> tg0_0:ctrl_ecc_readdataerror
	wire          hbm_0_example_design_ctrl_ecc_readdataerror_0_1_ctrl_ecc_readdataerror; // hbm_0_example_design:ctrl_ecc_readdataerror_0_1_ctrl_ecc_readdataerror -> tg0_1:ctrl_ecc_readdataerror
	wire          core_clk_iopll_locked_export;                                           // core_clk_iopll:locked -> hbm_0_example_design:ext_core_clk_locked
	wire          hbm_0_example_design_m2u_bridge_shiftwr;                                // hbm_0_example_design:shiftwr -> mem:shiftwr
	wire          hbm_0_example_design_m2u_bridge_updatewr;                               // hbm_0_example_design:updatewr -> mem:updatewr
	wire    [2:0] mem_m2u_bridge_temp;                                                    // mem:temp -> hbm_0_example_design:temp
	wire    [7:0] mem_m2u_bridge_wso;                                                     // mem:wso -> hbm_0_example_design:wso
	wire          mem_m2u_bridge_cattrip;                                                 // mem:cattrip -> hbm_0_example_design:cattrip
	wire          hbm_0_example_design_m2u_bridge_wrck;                                   // hbm_0_example_design:wrck -> mem:wrck
	wire          hbm_0_example_design_m2u_bridge_wrst_n;                                 // hbm_0_example_design:wrst_n -> mem:wrst_n
	wire          hbm_0_example_design_m2u_bridge_reset_n;                                // hbm_0_example_design:reset_n -> mem:reset_n
	wire          hbm_0_example_design_m2u_bridge_capturewr;                              // hbm_0_example_design:capturewr -> mem:capturewr
	wire          hbm_0_example_design_m2u_bridge_selectwir;                              // hbm_0_example_design:selectwir -> mem:selectwir
	wire          hbm_0_example_design_m2u_bridge_wsi;                                    // hbm_0_example_design:wsi -> mem:wsi
	wire    [3:0] hbm_0_example_design_mem_0_par;                                         // [] -> [hbm_0_example_design:par_0, mem:par_0]
	wire          hbm_0_example_design_mem_0_rr;                                          // hbm_0_example_design:rr_0 -> mem:rr_0
	wire          hbm_0_example_design_mem_0_ck_c;                                        // hbm_0_example_design:ck_c_0 -> mem:ck_c_0
	wire    [3:0] hbm_0_example_design_mem_0_wdqs_t;                                      // hbm_0_example_design:wdqs_t_0 -> mem:wdqs_t_0
	wire    [7:0] hbm_0_example_design_mem_0_c;                                           // hbm_0_example_design:c_0 -> mem:c_0
	wire    [3:0] mem_mem_0_rdqs_c;                                                       // mem:rdqs_c_0 -> hbm_0_example_design:rdqs_c_0
	wire   [15:0] hbm_0_example_design_mem_0_dm;                                          // [] -> [hbm_0_example_design:dm_0, mem:dm_0]
	wire          mem_mem_0_aerr;                                                         // mem:aerr_0 -> hbm_0_example_design:aerr_0
	wire   [15:0] hbm_0_example_design_mem_0_dbi;                                         // [] -> [hbm_0_example_design:dbi_0, mem:dbi_0]
	wire  [127:0] hbm_0_example_design_mem_0_dq;                                          // [] -> [hbm_0_example_design:dq_0, mem:dq_0]
	wire    [3:0] hbm_0_example_design_mem_0_derr;                                        // [] -> [hbm_0_example_design:derr_0, mem:derr_0]
	wire          hbm_0_example_design_mem_0_rc;                                          // hbm_0_example_design:rc_0 -> mem:rc_0
	wire    [5:0] hbm_0_example_design_mem_0_r;                                           // hbm_0_example_design:r_0 -> mem:r_0
	wire    [7:0] hbm_0_example_design_mem_0_rd;                                          // [] -> [hbm_0_example_design:rd_0, mem:rd_0]
	wire          hbm_0_example_design_mem_0_ck_t;                                        // hbm_0_example_design:ck_t_0 -> mem:ck_t_0
	wire    [3:0] hbm_0_example_design_mem_0_wdqs_c;                                      // hbm_0_example_design:wdqs_c_0 -> mem:wdqs_c_0
	wire    [3:0] mem_mem_0_rdqs_t;                                                       // mem:rdqs_t_0 -> hbm_0_example_design:rdqs_t_0
	wire          hbm_0_example_design_mem_0_cke;                                         // hbm_0_example_design:cke_0 -> mem:cke_0
	wire          reset_release_ip_ninit_done_ninit_done;                                 // reset_release_ip:ninit_done -> ninit_done_splitter:sig_input
	wire          ninit_done_splitter_sig_output_if_0_ninit_done;                         // ninit_done_splitter:sig_output_0 -> tg0_0:ninit_done
	wire          ninit_done_splitter_sig_output_if_1_ninit_done;                         // ninit_done_splitter:sig_output_1 -> tg0_1:ninit_done
	wire          hbm_0_example_design_status_local_cal_fail;                             // hbm_0_example_design:local_cal_fail -> sim_checker:local_cal_fail_0
	wire          hbm_0_example_design_status_local_cal_success;                          // hbm_0_example_design:local_cal_success -> sim_checker:local_cal_success_0
	wire          tg0_0_tg_status_traffic_gen_fail;                                       // tg0_0:traffic_gen_fail -> sim_checker:traffic_gen_fail_0
	wire          tg0_0_tg_status_traffic_gen_timeout;                                    // tg0_0:traffic_gen_timeout -> sim_checker:traffic_gen_timeout_0
	wire          tg0_0_tg_status_traffic_gen_pass;                                       // tg0_0:traffic_gen_pass -> sim_checker:traffic_gen_pass_0
	wire          tg0_1_tg_status_traffic_gen_fail;                                       // tg0_1:traffic_gen_fail -> sim_checker:traffic_gen_fail_1
	wire          tg0_1_tg_status_traffic_gen_timeout;                                    // tg0_1:traffic_gen_timeout -> sim_checker:traffic_gen_timeout_1
	wire          tg0_1_tg_status_traffic_gen_pass;                                       // tg0_1:traffic_gen_pass -> sim_checker:traffic_gen_pass_1
	wire          hbm_only_reset_source_reset_reset;                                      // hbm_only_reset_source:reset -> hbm_0_example_design:hbm_only_reset_in
	wire          global_reset_n_source_reset_reset;                                      // global_reset_n_source:reset -> [core_clk_iopll:rst, hbm_0_example_design:wmcrst_n_in]
	wire          hbm_0_example_design_wmcrst_n_0_reset;                                  // hbm_0_example_design:wmcrst_n_0_reset_n -> [tg0_0:wmcrst_n_in, tg0_1:wmcrst_n_in]

	ed_synth_core_clk_iopll core_clk_iopll (
		.refclk   (core_clk_source_clk_clk),            //   input,  width = 1,  refclk.clk
		.locked   (core_clk_iopll_locked_export),       //  output,  width = 1,  locked.export
		.rst      (~global_reset_n_source_reset_reset), //   input,  width = 1,   reset.reset
		.outclk_0 (core_clk_iopll_outclk0_clk)          //  output,  width = 1, outclk0.clk
	);

	ed_sim_core_clk_source core_clk_source (
		.clk (core_clk_source_clk_clk)  //  output,  width = 1, clk.clk
	);

	ed_sim_global_reset_n_source global_reset_n_source (
		.reset (global_reset_n_source_reset_reset), //  output,  width = 1, reset.reset_n
		.clk   (ref_clk_source_clk_clk)             //   input,  width = 1,   clk.clk
	);

	ed_synth_hbm_0_example_design hbm_0_example_design (
		.pll_ref_clk                                       (ref_clk_source_clk_clk),                                                 //   input,    width = 1,                pll_ref_clk.clk
		.ext_core_clk                                      (core_clk_iopll_outclk0_clk),                                             //   input,    width = 1,               ext_core_clk.clk
		.ext_core_clk_locked                               (core_clk_iopll_locked_export),                                           //   input,    width = 1,        ext_core_clk_locked.export
		.wmcrst_n_in                                       (global_reset_n_source_reset_reset),                                      //   input,    width = 1,                wmcrst_n_in.reset_n
		.hbm_only_reset_in                                 (hbm_only_reset_source_reset_reset),                                      //   input,    width = 1,          hbm_only_reset_in.reset
		.local_cal_success                                 (hbm_0_example_design_status_local_cal_success),                          //  output,    width = 1,                     status.local_cal_success
		.local_cal_fail                                    (hbm_0_example_design_status_local_cal_fail),                             //  output,    width = 1,                           .local_cal_fail
		.cal_lat                                           (),                                                                       //  output,    width = 3,                    cal_lat.cal_lat
		.ck_t_0                                            (hbm_0_example_design_mem_0_ck_t),                                        //  output,    width = 1,                      mem_0.ck_t
		.ck_c_0                                            (hbm_0_example_design_mem_0_ck_c),                                        //  output,    width = 1,                           .ck_c
		.cke_0                                             (hbm_0_example_design_mem_0_cke),                                         //  output,    width = 1,                           .cke
		.c_0                                               (hbm_0_example_design_mem_0_c),                                           //  output,    width = 8,                           .c
		.r_0                                               (hbm_0_example_design_mem_0_r),                                           //  output,    width = 6,                           .r
		.dq_0                                              (hbm_0_example_design_mem_0_dq),                                          //   inout,  width = 128,                           .dq
		.dm_0                                              (hbm_0_example_design_mem_0_dm),                                          //   inout,   width = 16,                           .dm
		.dbi_0                                             (hbm_0_example_design_mem_0_dbi),                                         //   inout,   width = 16,                           .dbi
		.par_0                                             (hbm_0_example_design_mem_0_par),                                         //   inout,    width = 4,                           .par
		.derr_0                                            (hbm_0_example_design_mem_0_derr),                                        //   inout,    width = 4,                           .derr
		.rdqs_t_0                                          (mem_mem_0_rdqs_t),                                                       //   input,    width = 4,                           .rdqs_t
		.rdqs_c_0                                          (mem_mem_0_rdqs_c),                                                       //   input,    width = 4,                           .rdqs_c
		.wdqs_t_0                                          (hbm_0_example_design_mem_0_wdqs_t),                                      //  output,    width = 4,                           .wdqs_t
		.wdqs_c_0                                          (hbm_0_example_design_mem_0_wdqs_c),                                      //  output,    width = 4,                           .wdqs_c
		.rd_0                                              (hbm_0_example_design_mem_0_rd),                                          //   inout,    width = 8,                           .rd
		.rr_0                                              (hbm_0_example_design_mem_0_rr),                                          //  output,    width = 1,                           .rr
		.rc_0                                              (hbm_0_example_design_mem_0_rc),                                          //  output,    width = 1,                           .rc
		.aerr_0                                            (mem_mem_0_aerr),                                                         //   input,    width = 1,                           .aerr
		.cattrip                                           (mem_m2u_bridge_cattrip),                                                 //   input,    width = 1,                 m2u_bridge.cattrip
		.temp                                              (mem_m2u_bridge_temp),                                                    //   input,    width = 3,                           .temp
		.wso                                               (mem_m2u_bridge_wso),                                                     //   input,    width = 8,                           .wso
		.reset_n                                           (hbm_0_example_design_m2u_bridge_reset_n),                                //  output,    width = 1,                           .reset_n
		.wrst_n                                            (hbm_0_example_design_m2u_bridge_wrst_n),                                 //  output,    width = 1,                           .wrst_n
		.wrck                                              (hbm_0_example_design_m2u_bridge_wrck),                                   //  output,    width = 1,                           .wrck
		.shiftwr                                           (hbm_0_example_design_m2u_bridge_shiftwr),                                //  output,    width = 1,                           .shiftwr
		.capturewr                                         (hbm_0_example_design_m2u_bridge_capturewr),                              //  output,    width = 1,                           .capturewr
		.updatewr                                          (hbm_0_example_design_m2u_bridge_updatewr),                               //  output,    width = 1,                           .updatewr
		.selectwir                                         (hbm_0_example_design_m2u_bridge_selectwir),                              //  output,    width = 1,                           .selectwir
		.wsi                                               (hbm_0_example_design_m2u_bridge_wsi),                                    //  output,    width = 1,                           .wsi
		.wmc_clk_0_clk                                     (hbm_0_example_design_wmc_clk_0_clk),                                     //  output,    width = 1,                  wmc_clk_0.clk
		.phy_clk_0_clk                                     (),                                                                       //  output,    width = 1,                  phy_clk_0.clk
		.wmcrst_n_0_reset_n                                (hbm_0_example_design_wmcrst_n_0_reset),                                  //  output,    width = 1,                 wmcrst_n_0.reset_n
		.ctrl_amm_0_1_waitrequest_n                        (tg0_1_ctrl_amm_waitrequest),                                             //  output,    width = 1,               ctrl_amm_0_1.waitrequest_n
		.ctrl_amm_0_1_read                                 (tg0_1_ctrl_amm_read),                                                    //   input,    width = 1,                           .read
		.ctrl_amm_0_1_write                                (tg0_1_ctrl_amm_write),                                                   //   input,    width = 1,                           .write
		.ctrl_amm_0_1_address                              (tg0_1_ctrl_amm_address),                                                 //   input,   width = 29,                           .address
		.ctrl_amm_0_1_readdata                             (tg0_1_ctrl_amm_readdata),                                                //  output,  width = 256,                           .readdata
		.ctrl_amm_0_1_writedata                            (tg0_1_ctrl_amm_writedata),                                               //   input,  width = 256,                           .writedata
		.ctrl_amm_0_1_burstcount                           (tg0_1_ctrl_amm_burstcount),                                              //   input,    width = 7,                           .burstcount
		.ctrl_amm_0_1_byteenable                           (tg0_1_ctrl_amm_byteenable),                                              //   input,   width = 32,                           .byteenable
		.ctrl_amm_0_1_readdatavalid                        (tg0_1_ctrl_amm_readdatavalid),                                           //  output,    width = 1,                           .readdatavalid
		.ctrl_amm_0_0_waitrequest_n                        (tg0_0_ctrl_amm_waitrequest),                                             //  output,    width = 1,               ctrl_amm_0_0.waitrequest_n
		.ctrl_amm_0_0_read                                 (tg0_0_ctrl_amm_read),                                                    //   input,    width = 1,                           .read
		.ctrl_amm_0_0_write                                (tg0_0_ctrl_amm_write),                                                   //   input,    width = 1,                           .write
		.ctrl_amm_0_0_address                              (tg0_0_ctrl_amm_address),                                                 //   input,   width = 29,                           .address
		.ctrl_amm_0_0_readdata                             (tg0_0_ctrl_amm_readdata),                                                //  output,  width = 256,                           .readdata
		.ctrl_amm_0_0_writedata                            (tg0_0_ctrl_amm_writedata),                                               //   input,  width = 256,                           .writedata
		.ctrl_amm_0_0_burstcount                           (tg0_0_ctrl_amm_burstcount),                                              //   input,    width = 7,                           .burstcount
		.ctrl_amm_0_0_byteenable                           (tg0_0_ctrl_amm_byteenable),                                              //   input,   width = 32,                           .byteenable
		.ctrl_amm_0_0_readdatavalid                        (tg0_0_ctrl_amm_readdatavalid),                                           //  output,    width = 1,                           .readdatavalid
		.ctrl_ecc_readdataerror_0_1_ctrl_ecc_readdataerror (hbm_0_example_design_ctrl_ecc_readdataerror_0_1_ctrl_ecc_readdataerror), //  output,    width = 1, ctrl_ecc_readdataerror_0_1.ctrl_ecc_readdataerror
		.ctrl_ecc_readdataerror_0_0_ctrl_ecc_readdataerror (hbm_0_example_design_ctrl_ecc_readdataerror_0_0_ctrl_ecc_readdataerror), //  output,    width = 1, ctrl_ecc_readdataerror_0_0.ctrl_ecc_readdataerror
		.apb_0_ur_paddr                                    (tg0_0_apb_ur_paddr),                                                     //   input,   width = 16,                      apb_0.ur_paddr
		.apb_0_ur_psel                                     (tg0_0_apb_ur_psel),                                                      //   input,    width = 1,                           .ur_psel
		.apb_0_ur_penable                                  (tg0_0_apb_ur_penable),                                                   //   input,    width = 1,                           .ur_penable
		.apb_0_ur_pwrite                                   (tg0_0_apb_ur_pwrite),                                                    //   input,    width = 1,                           .ur_pwrite
		.apb_0_ur_pwdata                                   (tg0_0_apb_ur_pwdata),                                                    //   input,   width = 16,                           .ur_pwdata
		.apb_0_ur_pstrb                                    (tg0_0_apb_ur_pstrb),                                                     //   input,    width = 2,                           .ur_pstrb
		.apb_0_ur_prready                                  (hbm_0_example_design_apb_0_ur_prready),                                  //  output,    width = 1,                           .ur_prready
		.apb_0_ur_prdata                                   (hbm_0_example_design_apb_0_ur_prdata)                                    //  output,   width = 16,                           .ur_prdata
	);

	ed_sim_hbm_only_reset_source hbm_only_reset_source (
		.reset (hbm_only_reset_source_reset_reset), //  output,  width = 1, reset.reset
		.clk   (ref_clk_source_clk_clk)             //   input,  width = 1,   clk.clk
	);

	ed_sim_mem mem (
		.ck_t_0    (hbm_0_example_design_mem_0_ck_t),           //   input,    width = 1,      mem_0.ck_t
		.ck_c_0    (hbm_0_example_design_mem_0_ck_c),           //   input,    width = 1,           .ck_c
		.cke_0     (hbm_0_example_design_mem_0_cke),            //   input,    width = 1,           .cke
		.c_0       (hbm_0_example_design_mem_0_c),              //   input,    width = 8,           .c
		.r_0       (hbm_0_example_design_mem_0_r),              //   input,    width = 6,           .r
		.dq_0      (hbm_0_example_design_mem_0_dq),             //   inout,  width = 128,           .dq
		.dm_0      (hbm_0_example_design_mem_0_dm),             //   inout,   width = 16,           .dm
		.dbi_0     (hbm_0_example_design_mem_0_dbi),            //   inout,   width = 16,           .dbi
		.par_0     (hbm_0_example_design_mem_0_par),            //   inout,    width = 4,           .par
		.derr_0    (hbm_0_example_design_mem_0_derr),           //   inout,    width = 4,           .derr
		.rdqs_t_0  (mem_mem_0_rdqs_t),                          //  output,    width = 4,           .rdqs_t
		.rdqs_c_0  (mem_mem_0_rdqs_c),                          //  output,    width = 4,           .rdqs_c
		.wdqs_t_0  (hbm_0_example_design_mem_0_wdqs_t),         //   input,    width = 4,           .wdqs_t
		.wdqs_c_0  (hbm_0_example_design_mem_0_wdqs_c),         //   input,    width = 4,           .wdqs_c
		.rd_0      (hbm_0_example_design_mem_0_rd),             //   inout,    width = 8,           .rd
		.rr_0      (hbm_0_example_design_mem_0_rr),             //   input,    width = 1,           .rr
		.rc_0      (hbm_0_example_design_mem_0_rc),             //   input,    width = 1,           .rc
		.aerr_0    (mem_mem_0_aerr),                            //  output,    width = 1,           .aerr
		.cattrip   (mem_m2u_bridge_cattrip),                    //  output,    width = 1, m2u_bridge.cattrip
		.temp      (mem_m2u_bridge_temp),                       //  output,    width = 3,           .temp
		.wso       (mem_m2u_bridge_wso),                        //  output,    width = 8,           .wso
		.reset_n   (hbm_0_example_design_m2u_bridge_reset_n),   //   input,    width = 1,           .reset_n
		.wrst_n    (hbm_0_example_design_m2u_bridge_wrst_n),    //   input,    width = 1,           .wrst_n
		.wrck      (hbm_0_example_design_m2u_bridge_wrck),      //   input,    width = 1,           .wrck
		.shiftwr   (hbm_0_example_design_m2u_bridge_shiftwr),   //   input,    width = 1,           .shiftwr
		.capturewr (hbm_0_example_design_m2u_bridge_capturewr), //   input,    width = 1,           .capturewr
		.updatewr  (hbm_0_example_design_m2u_bridge_updatewr),  //   input,    width = 1,           .updatewr
		.selectwir (hbm_0_example_design_m2u_bridge_selectwir), //   input,    width = 1,           .selectwir
		.wsi       (hbm_0_example_design_m2u_bridge_wsi)        //   input,    width = 1,           .wsi
	);

	ed_synth_ninit_done_splitter ninit_done_splitter (
		.sig_input    (reset_release_ip_ninit_done_ninit_done),         //   input,  width = 1,    sig_input_if.ninit_done
		.sig_output_0 (ninit_done_splitter_sig_output_if_0_ninit_done), //  output,  width = 1, sig_output_if_0.ninit_done
		.sig_output_1 (ninit_done_splitter_sig_output_if_1_ninit_done)  //  output,  width = 1, sig_output_if_1.ninit_done
	);

	ed_sim_ref_clk_source ref_clk_source (
		.clk (ref_clk_source_clk_clk)  //  output,  width = 1, clk.clk
	);

	ed_synth_reset_release_ip reset_release_ip (
		.ninit_done (reset_release_ip_ninit_done_ninit_done)  //  output,  width = 1, ninit_done.ninit_done
	);

	ed_sim_sim_checker sim_checker (
		.traffic_gen_pass_0    (tg0_0_tg_status_traffic_gen_pass),              //   input,  width = 1, tg_status_0.traffic_gen_pass
		.traffic_gen_fail_0    (tg0_0_tg_status_traffic_gen_fail),              //   input,  width = 1,            .traffic_gen_fail
		.traffic_gen_timeout_0 (tg0_0_tg_status_traffic_gen_timeout),           //   input,  width = 1,            .traffic_gen_timeout
		.traffic_gen_pass_1    (tg0_1_tg_status_traffic_gen_pass),              //   input,  width = 1, tg_status_1.traffic_gen_pass
		.traffic_gen_fail_1    (tg0_1_tg_status_traffic_gen_fail),              //   input,  width = 1,            .traffic_gen_fail
		.traffic_gen_timeout_1 (tg0_1_tg_status_traffic_gen_timeout),           //   input,  width = 1,            .traffic_gen_timeout
		.traffic_gen_pass      (sim_checker_traffic_gen_pass),                  //  output,  width = 1,   tg_status.traffic_gen_pass
		.traffic_gen_fail      (sim_checker_traffic_gen_fail),                  //  output,  width = 1,            .traffic_gen_fail
		.traffic_gen_timeout   (sim_checker_traffic_gen_timeout),               //  output,  width = 1,            .traffic_gen_timeout
		.local_cal_success_0   (hbm_0_example_design_status_local_cal_success), //   input,  width = 1,    status_0.local_cal_success
		.local_cal_fail_0      (hbm_0_example_design_status_local_cal_fail),    //   input,  width = 1,            .local_cal_fail
		.local_cal_success     (cal_status_checker_local_cal_success),          //  output,  width = 1,      status.local_cal_success
		.local_cal_fail        (cal_status_checker_local_cal_fail)              //  output,  width = 1,            .local_cal_fail
	);

	ed_synth_tg0_0 tg0_0 (
		.ninit_done             (ninit_done_splitter_sig_output_if_0_ninit_done),                         //   input,    width = 1,             ninit_done.ninit_done
		.wmc_clk_in             (hbm_0_example_design_wmc_clk_0_clk),                                     //   input,    width = 1,             wmc_clk_in.clk
		.wmcrst_n_in            (hbm_0_example_design_wmcrst_n_0_reset),                                  //   input,    width = 1,            wmcrst_n_in.reset_n
		.amm_ready              (tg0_0_ctrl_amm_waitrequest),                                             //   input,    width = 1,               ctrl_amm.waitrequest_n
		.amm_read               (tg0_0_ctrl_amm_read),                                                    //  output,    width = 1,                       .read
		.amm_write              (tg0_0_ctrl_amm_write),                                                   //  output,    width = 1,                       .write
		.amm_address            (tg0_0_ctrl_amm_address),                                                 //  output,   width = 29,                       .address
		.amm_readdata           (tg0_0_ctrl_amm_readdata),                                                //   input,  width = 256,                       .readdata
		.amm_writedata          (tg0_0_ctrl_amm_writedata),                                               //  output,  width = 256,                       .writedata
		.amm_burstcount         (tg0_0_ctrl_amm_burstcount),                                              //  output,    width = 7,                       .burstcount
		.amm_byteenable         (tg0_0_ctrl_amm_byteenable),                                              //  output,   width = 32,                       .byteenable
		.amm_readdatavalid      (tg0_0_ctrl_amm_readdatavalid),                                           //   input,    width = 1,                       .readdatavalid
		.traffic_gen_pass       (tg0_0_tg_status_traffic_gen_pass),                                       //  output,    width = 1,              tg_status.traffic_gen_pass
		.traffic_gen_fail       (tg0_0_tg_status_traffic_gen_fail),                                       //  output,    width = 1,                       .traffic_gen_fail
		.traffic_gen_timeout    (tg0_0_tg_status_traffic_gen_timeout),                                    //  output,    width = 1,                       .traffic_gen_timeout
		.ctrl_ecc_readdataerror (hbm_0_example_design_ctrl_ecc_readdataerror_0_0_ctrl_ecc_readdataerror), //   input,    width = 1, ctrl_ecc_readdataerror.ctrl_ecc_readdataerror
		.ur_paddr               (tg0_0_apb_ur_paddr),                                                     //  output,   width = 16,                    apb.ur_paddr
		.ur_psel                (tg0_0_apb_ur_psel),                                                      //  output,    width = 1,                       .ur_psel
		.ur_penable             (tg0_0_apb_ur_penable),                                                   //  output,    width = 1,                       .ur_penable
		.ur_pwrite              (tg0_0_apb_ur_pwrite),                                                    //  output,    width = 1,                       .ur_pwrite
		.ur_pwdata              (tg0_0_apb_ur_pwdata),                                                    //  output,   width = 16,                       .ur_pwdata
		.ur_pstrb               (tg0_0_apb_ur_pstrb),                                                     //  output,    width = 2,                       .ur_pstrb
		.ur_prready             (hbm_0_example_design_apb_0_ur_prready),                                  //   input,    width = 1,                       .ur_prready
		.ur_prdata              (hbm_0_example_design_apb_0_ur_prdata)                                    //   input,   width = 16,                       .ur_prdata
	);

	ed_synth_tg0_1 tg0_1 (
		.ninit_done             (ninit_done_splitter_sig_output_if_1_ninit_done),                         //   input,    width = 1,             ninit_done.ninit_done
		.wmc_clk_in             (hbm_0_example_design_wmc_clk_0_clk),                                     //   input,    width = 1,             wmc_clk_in.clk
		.wmcrst_n_in            (hbm_0_example_design_wmcrst_n_0_reset),                                  //   input,    width = 1,            wmcrst_n_in.reset_n
		.amm_ready              (tg0_1_ctrl_amm_waitrequest),                                             //   input,    width = 1,               ctrl_amm.waitrequest_n
		.amm_read               (tg0_1_ctrl_amm_read),                                                    //  output,    width = 1,                       .read
		.amm_write              (tg0_1_ctrl_amm_write),                                                   //  output,    width = 1,                       .write
		.amm_address            (tg0_1_ctrl_amm_address),                                                 //  output,   width = 29,                       .address
		.amm_readdata           (tg0_1_ctrl_amm_readdata),                                                //   input,  width = 256,                       .readdata
		.amm_writedata          (tg0_1_ctrl_amm_writedata),                                               //  output,  width = 256,                       .writedata
		.amm_burstcount         (tg0_1_ctrl_amm_burstcount),                                              //  output,    width = 7,                       .burstcount
		.amm_byteenable         (tg0_1_ctrl_amm_byteenable),                                              //  output,   width = 32,                       .byteenable
		.amm_readdatavalid      (tg0_1_ctrl_amm_readdatavalid),                                           //   input,    width = 1,                       .readdatavalid
		.traffic_gen_pass       (tg0_1_tg_status_traffic_gen_pass),                                       //  output,    width = 1,              tg_status.traffic_gen_pass
		.traffic_gen_fail       (tg0_1_tg_status_traffic_gen_fail),                                       //  output,    width = 1,                       .traffic_gen_fail
		.traffic_gen_timeout    (tg0_1_tg_status_traffic_gen_timeout),                                    //  output,    width = 1,                       .traffic_gen_timeout
		.ctrl_ecc_readdataerror (hbm_0_example_design_ctrl_ecc_readdataerror_0_1_ctrl_ecc_readdataerror)  //   input,    width = 1, ctrl_ecc_readdataerror.ctrl_ecc_readdataerror
	);

endmodule
